library verilog;
use verilog.vl_types.all;
entity topmodule_nios2_vlg_vec_tst is
end topmodule_nios2_vlg_vec_tst;
