library verilog;
use verilog.vl_types.all;
entity IP_wrapper_vlg_vec_tst is
end IP_wrapper_vlg_vec_tst;
