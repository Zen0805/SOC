
module message_scheduler (
    input wire          clk,
    input wire          reset_n,         // Reset tích cực thấp
    input wire          start_new_block, // Báo hiệu bắt đầu block mới
    input wire [5:0]    round_t,         // Vòng lặp hiện tại (0-63)
    input wire [31:0]   message_word_in, // Dữ liệu M[i] để load
    input wire [3:0]    message_word_addr,// Địa chỉ (0-15) của M[i] đang load
    input wire          write_enable_in, // Cho phép ghi message_word_in vào memory
    output wire [31:0]  Wt_out           // W[t] tương ứng với round_t
);

    // --- Internal Signals ---
    reg [31:0] W_memory [15:0];     // Bộ nhớ lưu 16 từ W[t-16] đến W[t-1]
    reg [31:0] reg_w;               // Lưu kết quả cộng trung gian và W[t] cuối cùng
    reg [1:0] calc_cycle;           // 0: s1, 1: s2, 2: s3, 3: s4
    reg calculation_active;         // Đánh dấu đang tính toán 4 chu kỳ
    reg [31:0] prev_wt;             // Lưu W[t] của vòng trước để ghi ở vòng sau

    wire [31:0] mem_out_t_minus_16;
    wire [31:0] mem_out_t_minus_15;
    wire [31:0] mem_out_t_minus_7;
    wire [31:0] mem_out_t_minus_2;

    wire [3:0] addr_t_minus_16;
    wire [3:0] addr_t_minus_15;
    wire [3:0] addr_t_minus_7;
    wire [3:0] addr_t_minus_2;
    wire [3:0] write_addr;

    wire [31:0] sigma0_result;
    wire [31:0] sigma1_result;

    wire [31:0] adder_in_a;         // Đầu vào A của bộ cộng
    wire [31:0] adder_in_b;         // Đầu vào B của bộ cộng
    wire [31:0] adder_sum_out;      // Kết quả từ bộ cộng

    // --- Tính toán địa chỉ Memory (Modulo 16) ---
    assign addr_t_minus_16 = round_t[3:0];           // W[t-16] = t mod 16
    assign addr_t_minus_15 = (round_t - 6'd15) & 4'hF;// (t-15) mod 16
    assign addr_t_minus_7  = (round_t - 6'd7) & 4'hF; // (t-7) mod 16
    assign addr_t_minus_2  = (round_t - 6'd2) & 4'hF; // (t-2) mod 16
    assign write_addr      = addr_t_minus_16;        // Ghi đè lên W[t-16]

    // --- Đọc dữ liệu từ Memory ---
    assign mem_out_t_minus_16 = W_memory[addr_t_minus_16];
    assign mem_out_t_minus_15 = W_memory[addr_t_minus_15];
    assign mem_out_t_minus_7  = W_memory[addr_t_minus_7];
    assign mem_out_t_minus_2  = W_memory[addr_t_minus_2];

    // --- Khởi tạo các hàm Sigma ---
    sigma0_func_schedule u_sigma0 (.x(mem_out_t_minus_15), .out(sigma0_result));
    sigma1_func_schedule u_sigma1 (.x(mem_out_t_minus_2),  .out(sigma1_result));

    // --- Khởi tạo bộ cộng 32-bit ---
    adder_32bit u_adder (.a(adder_in_a), .b(adder_in_b), .sum(adder_sum_out));

    // --- Logic chọn đầu vào cho bộ cộng (Combinational) ---
    assign adder_in_a = (calculation_active && calc_cycle == 2'b00) ? mem_out_t_minus_16 :
                        (calculation_active && (calc_cycle == 2'b01 || calc_cycle == 2'b10)) ? reg_w :
                        32'b0;

    assign adder_in_b = (calculation_active && calc_cycle == 2'b00) ? sigma0_result :
                        (calculation_active && calc_cycle == 2'b01) ? mem_out_t_minus_7 :
                        (calculation_active && calc_cycle == 2'b10) ? sigma1_result :
                        32'b0;

    // --- Logic điều khiển và cập nhật trạng thái (Sequential) ---
    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            calc_cycle <= 2'b00;
            reg_w <= 32'b0;
            calculation_active <= 1'b0;
            prev_wt <= 32'b0;
        end else begin
            // --- Ghi dữ liệu đầu vào (M[i]) vào memory ---
            if (write_enable_in) begin
                W_memory[message_word_addr] <= message_word_in;
            end

            // --- Tính toán W[t] cho t >= 16 ---
            if (round_t >= 6'd16) begin
                if (!calculation_active) begin // Bắt đầu tính toán cho round mới
                    calculation_active <= 1'b1;
                    calc_cycle <= 2'b00;
                    // Ghi W[t-1] từ vòng trước vào bộ nhớ ở cycle 0 của vòng mới
                    if (round_t > 6'd16) begin
                        W_memory[write_addr] <= prev_wt;
                        $display("[%0t] Writing W[%0d] = 0x%h to memory at addr %0d", $time, round_t - 1, prev_wt, write_addr);
                    end
                end else begin // Đang trong quá trình tính toán
                    if (calc_cycle == 2'b00 || calc_cycle == 2'b01 || calc_cycle == 2'b10) begin
                        reg_w <= adder_sum_out;
                    end
                    case (calc_cycle)
                        2'b00: begin
                            calc_cycle <= 2'b01;
                            $display("[%0t] Calculating W[%0d]:", $time, round_t);
                            $display("  W[t-16] = 0x%h", mem_out_t_minus_16);
                            $display("  W[t-15] = 0x%h", mem_out_t_minus_15);
                            $display("  W[t-7]  = 0x%h", mem_out_t_minus_7);
                            $display("  W[t-2]  = 0x%h", mem_out_t_minus_2);
                            $display("  σ0(W[t-15]) = 0x%h", sigma0_result);
                            $display("  σ1(W[t-2])  = 0x%h", sigma1_result);
                        end
                        2'b01: calc_cycle <= 2'b10;
                        2'b10: begin
                            calc_cycle <= 2'b11;
                            prev_wt <= adder_sum_out; // Lưu W[t] cho lần ghi tiếp theo
                        end
                        2'b11: begin
                            calc_cycle <= 2'b00;
                            calculation_active <= 1'b0;
                        end
                        default: begin
                            calc_cycle <= 2'b00;
                            calculation_active <= 1'b0;
                        end
                    endcase
                end
            end else begin // round_t < 16
                calculation_active <= 1'b0;
                calc_cycle <= 2'b00;
            end
        end
    end

    // --- Logic chọn đầu ra Wt_out (Combinational) ---
    assign Wt_out = (round_t < 6'd16) ? W_memory[addr_t_minus_16] : reg_w;

endmodule

