library verilog;
use verilog.vl_types.all;
entity sha256_optimizePowerAreaVerilog_vlg_vec_tst is
end sha256_optimizePowerAreaVerilog_vlg_vec_tst;
