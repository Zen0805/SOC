//-----------------------------------------------------------------------------
// Module: Sigma1_func_for_compression
// Chức năng: Tính hàm Sigma1 hoa (Σ₁) của SHA-256 (dùng trong compression).
//            Σ₁(x) = ROTR⁶(x) ^ ROTR¹¹(x) ^ ROTR²⁵(x)
//-----------------------------------------------------------------------------
module sigma1_func_compression (
    input wire [31:0] x,
    output wire [31:0] out
);

    wire [31:0] rotr6_x;
    wire [31:0] rotr11_x;
    wire [31:0] rotr25_x;

    // Rotate Right 6 bits: {lower 6 bits, upper 26 bits}
    assign rotr6_x  = {x[5:0], x[31:6]};
    // Rotate Right 11 bits: {lower 11 bits, upper 21 bits}
    assign rotr11_x = {x[10:0], x[31:11]};
    // Rotate Right 25 bits: {lower 25 bits, upper 7 bits}
    assign rotr25_x = {x[24:0], x[31:25]};

    // XOR các kết quả lại
    assign out = rotr6_x ^ rotr11_x ^ rotr25_x;

endmodule